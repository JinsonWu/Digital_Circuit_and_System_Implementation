module Lab01(
  // Input signals
  in_number1,
  in_number2,
  in_number3,
  in_number4,
  // Output signals
  out_number1,
  out_number2
);

//---------------------------------------------------------------------
//   INPUT AND OUTPUT DECLARATION                         
//---------------------------------------------------------------------
input [3:0] in_number1,in_number2,in_number3,in_number4;

output logic [4:0] out_number1,out_number2;


endmodule
